
module test_probe (
	source,
	probe,
	source_clk);	

	output	[86:0]	source;
	input	[85:0]	probe;
	input		source_clk;
endmodule
